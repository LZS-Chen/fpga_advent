/**
 * Step 1: Blinker
 * DONE
 */

`default_nettype none

module SOC (
    input  CLK,        // system clock 
    input  RESET,      // reset button
   //  output LED // system LEDs
    output [4:0] LEDS, // system LEDs

    input  RXD,        // UART receive
    output TXD         // UART transmit
);


// A blinker that counts on 5 bits, wired to the 5 LEDs
   reg [4:0] count = 0;
   always @(posedge CLK) begin
      count <= count + 1;
   end
   assign LEDS = count;
   assign TXD  = 1'b0; // not used for now
endmodule
